// Wrapper for vivado_system. This matches the signals' names in XPS with
// those of Vivado.

module system (
  inout [53:0] processing_system7_0_MIO,
  input processing_system7_0_PS_SRSTB,
  input processing_system7_0_PS_CLK,
  input processing_system7_0_PS_PORB,
  inout processing_system7_0_DDR_Clk,
  inout processing_system7_0_DDR_Clk_n,
  inout processing_system7_0_DDR_CKE,
  inout processing_system7_0_DDR_CS_n,
  inout processing_system7_0_DDR_RAS_n,
  inout processing_system7_0_DDR_CAS_n,
  output processing_system7_0_DDR_WEB,
  inout [2:0] processing_system7_0_DDR_BankAddr,
  inout [14:0] processing_system7_0_DDR_Addr,
  inout processing_system7_0_DDR_ODT,
  inout processing_system7_0_DDR_DRSTB,
  inout [31:0] processing_system7_0_DDR_DQ,
  inout [3:0] processing_system7_0_DDR_DM,
  inout [3:0] processing_system7_0_DDR_DQS,
  inout [3:0] processing_system7_0_DDR_DQS_n,
  inout processing_system7_0_DDR_VRN,
  inout processing_system7_0_DDR_VRP,
 /* output xillybus_bus_clk,
  output xillybus_bus_rst_n,
  output [31:0] xillybus_S_AXI_AWADDR,
  output xillybus_S_AXI_AWVALID,
  output [31:0] xillybus_S_AXI_WDATA,
  output [3:0] xillybus_S_AXI_WSTRB,
  output xillybus_S_AXI_WVALID,
  output xillybus_S_AXI_BREADY,
  output [31:0] xillybus_S_AXI_ARADDR,
  output xillybus_S_AXI_ARVALID,
  output xillybus_S_AXI_RREADY,
  input xillybus_S_AXI_ARREADY,
  input [31:0] xillybus_S_AXI_RDATA,
  input [1:0] xillybus_S_AXI_RRESP,
  input xillybus_S_AXI_RVALID,
  input xillybus_S_AXI_WREADY,
  input [1:0] xillybus_S_AXI_BRESP,
  input xillybus_S_AXI_BVALID,
  input xillybus_S_AXI_AWREADY,
  output xillybus_M_AXI_ARREADY,
  input xillybus_M_AXI_ARVALID,
  input [31:0] xillybus_M_AXI_ARADDR,
  input [3:0] xillybus_M_AXI_ARLEN,
  input [2:0] xillybus_M_AXI_ARSIZE,
  input [1:0] xillybus_M_AXI_ARBURST,
  input [2:0] xillybus_M_AXI_ARPROT,
  input [3:0] xillybus_M_AXI_ARCACHE,
  input xillybus_M_AXI_RREADY,
  output xillybus_M_AXI_RVALID,
  output [63:0] xillybus_M_AXI_RDATA,
  output [1:0] xillybus_M_AXI_RRESP,
  output xillybus_M_AXI_RLAST,
  output xillybus_M_AXI_AWREADY,
  input xillybus_M_AXI_AWVALID,
  input [31:0] xillybus_M_AXI_AWADDR,
  input [3:0] xillybus_M_AXI_AWLEN,
  input [2:0] xillybus_M_AXI_AWSIZE,
  input [1:0] xillybus_M_AXI_AWBURST,
  input [2:0] xillybus_M_AXI_AWPROT,
  input [3:0] xillybus_M_AXI_AWCACHE,
  output xillybus_M_AXI_WREADY,
  input xillybus_M_AXI_WVALID,
  input [63:0] xillybus_M_AXI_WDATA,
  input [7:0] xillybus_M_AXI_WSTRB,
  input xillybus_M_AXI_WLAST,
  input xillybus_M_AXI_BREADY,
  output xillybus_M_AXI_BVALID,
  output [1:0] xillybus_M_AXI_BRESP,
  input xillybus_host_interrupt, */
  inout [55:0] processing_system7_0_GPIO,
  input processing_system7_0_USB0_VBUS_PWRFAULT,
  output xillybus_lite_0_user_clk_pin,
  output xillybus_lite_0_user_wren_pin,
  output [3:0] xillybus_lite_0_user_wstrb_pin,
  output xillybus_lite_0_user_rden_pin,
  input [31:0] xillybus_lite_0_user_rd_data_pin,
  output [31:0] xillybus_lite_0_user_wr_data_pin,
  output [31:0] xillybus_lite_0_user_addr_pin,
  input xillybus_lite_0_user_irq_pin, 
  
  output mdio_phy_mdc,
  inout mdio_phy_io,
  output [1:0] rmii2phy_txd,
  output rmii2phy_tx_en,
  input phy2rmii_rx_er,
  input phy2rmii_crs_dv,
  input [1:0] phy2rmii_rxd,
  input ethclk50,
  input reset_rtl,
  
  output [5:0] testmii
  
);
wire mdio_phy_o, mdio_phy_i, mdio_phy_t; 
     assign testmii[2] = mdio_phy_mdc;
     assign testmii[3] = mdio_phy_i;
     assign testmii[4] = mdio_phy_o;
     assign testmii[5] = mdio_phy_t;
/*
       wire mdio_phy_o, mdio_phy_i, mdio_phy_t; 
	   assign mdio_phy_i = mdio_phy_io; 
	   assign mdio_phy_io = mdio_phy_t ? 1'bz :  mdio_phy_o;
*/
   wire [55:0] gpio_tri_i, gpio_tri_o, gpio_tri_t;
   genvar      i;

   generate
      for (i=0; i<56; i=i+1)
	begin: gpio
	   assign gpio_tri_i[i] = processing_system7_0_GPIO[i]; 
	   assign processing_system7_0_GPIO[i] = gpio_tri_t[i] ? 1'bz :
						 gpio_tri_o[i];
	end
   endgenerate
   
     IOBUF mdio_rtl_mdio_iobuf
        (.I(mdio_phy_o),
         .IO(mdio_phy_io),
         .O(mdio_phy_i),
         .T(mdio_phy_t));
   
vivado_system vivado_system_i
       (.DDR_addr(processing_system7_0_DDR_Addr),
        .DDR_ba(processing_system7_0_DDR_BankAddr),
        .DDR_cas_n(processing_system7_0_DDR_CAS_n),
        .DDR_ck_n(processing_system7_0_DDR_Clk_n),
        .DDR_ck_p(processing_system7_0_DDR_Clk_p),
        .DDR_cke(processing_system7_0_DDR_CKE),
        .DDR_cs_n(processing_system7_0_DDR_CS_n),
        .DDR_dm(processing_system7_0_DDR_DM),
        .DDR_dq(processing_system7_0_DDR_DQ),
        .DDR_dqs_n(processing_system7_0_DDR_DQS_n),
        .DDR_dqs_p(processing_system7_0_DDR_DQS),
        .DDR_odt(processing_system7_0_DDR_ODT),
        .DDR_ras_n(processing_system7_0_DDR_RAS_n),
        .DDR_reset_n(processing_system7_0_DDR_DRSTB),
        .DDR_we_n(processing_system7_0_DDR_WEB),
        .FIXED_IO_ddr_vrn(processing_system7_0_DDR_VRN),
        .FIXED_IO_ddr_vrp(processing_system7_0_DDR_VRP),
        .FIXED_IO_mio(processing_system7_0_MIO),
        .FIXED_IO_ps_clk(processing_system7_0_PS_CLK),
        .FIXED_IO_ps_porb(processing_system7_0_PS_PORB),
        .FIXED_IO_ps_srstb(processing_system7_0_PS_SRSTB),
        .GPIO_0_tri_i(gpio_tri_i),
        .GPIO_0_tri_o(gpio_tri_o),
        .GPIO_0_tri_t(gpio_tri_t),
        .USBIND_0_port_indctl(),
        .USBIND_0_vbus_pwrfault(processing_system7_0_USB0_VBUS_PWRFAULT),
        .USBIND_0_vbus_pwrselect(),
        .user_addr(xillybus_lite_0_user_addr_pin),
        .user_clk(xillybus_lite_0_user_clk_pin),
        .user_irq(xillybus_lite_0_user_irq_pin),
        .user_rd_data(xillybus_lite_0_user_rd_data_pin),
        .user_rden(xillybus_lite_0_user_rden_pin),
        .user_wr_data(xillybus_lite_0_user_wr_data_pin),
        .user_wren(xillybus_lite_0_user_wren_pin),
        .user_wstrb(xillybus_lite_0_user_wstrb_pin),
  /*      .xillybus_M_AXI_araddr(xillybus_M_AXI_ARADDR),
        .xillybus_M_AXI_arburst(xillybus_M_AXI_ARBURST),
        .xillybus_M_AXI_arcache(xillybus_M_AXI_ARCACHE),
        .xillybus_M_AXI_arlen(xillybus_M_AXI_ARLEN),
        .xillybus_M_AXI_arprot(xillybus_M_AXI_ARPROT),
        .xillybus_M_AXI_arready(xillybus_M_AXI_ARREADY),
        .xillybus_M_AXI_arsize(xillybus_M_AXI_ARSIZE),
        .xillybus_M_AXI_arvalid(xillybus_M_AXI_ARVALID),
        .xillybus_M_AXI_awaddr(xillybus_M_AXI_AWADDR),
        .xillybus_M_AXI_awburst(xillybus_M_AXI_AWBURST),
        .xillybus_M_AXI_awcache(xillybus_M_AXI_AWCACHE),
        .xillybus_M_AXI_awlen(xillybus_M_AXI_AWLEN),
        .xillybus_M_AXI_awprot(xillybus_M_AXI_AWPROT),
        .xillybus_M_AXI_awready(xillybus_M_AXI_AWREADY),
        .xillybus_M_AXI_awsize(xillybus_M_AXI_AWSIZE),
        .xillybus_M_AXI_awvalid(xillybus_M_AXI_AWVALID),
        .xillybus_M_AXI_bready(xillybus_M_AXI_BREADY),
        .xillybus_M_AXI_bresp(xillybus_M_AXI_BRESP),
        .xillybus_M_AXI_bvalid(xillybus_M_AXI_BVALID),
        .xillybus_M_AXI_rdata(xillybus_M_AXI_RDATA),
        .xillybus_M_AXI_rlast(xillybus_M_AXI_RLAST),
        .xillybus_M_AXI_rready(xillybus_M_AXI_RREADY),
        .xillybus_M_AXI_rresp(xillybus_M_AXI_RRESP),
        .xillybus_M_AXI_rvalid(xillybus_M_AXI_RVALID),
        .xillybus_M_AXI_wdata(xillybus_M_AXI_WDATA),
        .xillybus_M_AXI_wlast(xillybus_M_AXI_WLAST),
        .xillybus_M_AXI_wready(xillybus_M_AXI_WREADY),
        .xillybus_M_AXI_wstrb(xillybus_M_AXI_WSTRB),
        .xillybus_M_AXI_wvalid(xillybus_M_AXI_WVALID),
        .xillybus_S_AXI_araddr(xillybus_S_AXI_ARADDR),
        .xillybus_S_AXI_arready(xillybus_S_AXI_ARREADY),
        .xillybus_S_AXI_arvalid(xillybus_S_AXI_ARVALID),
        .xillybus_S_AXI_awaddr(xillybus_S_AXI_AWADDR),
        .xillybus_S_AXI_awready(xillybus_S_AXI_AWREADY),
        .xillybus_S_AXI_awvalid(xillybus_S_AXI_AWVALID),
        .xillybus_S_AXI_bready(xillybus_S_AXI_BREADY),
        .xillybus_S_AXI_bresp(xillybus_S_AXI_BRESP),
        .xillybus_S_AXI_bvalid(xillybus_S_AXI_BVALID),
        .xillybus_S_AXI_rdata(xillybus_S_AXI_RDATA),
        .xillybus_S_AXI_rready(xillybus_S_AXI_RREADY),
        .xillybus_S_AXI_rresp(xillybus_S_AXI_RRESP),
        .xillybus_S_AXI_rvalid(xillybus_S_AXI_RVALID),
        .xillybus_S_AXI_wdata(xillybus_S_AXI_WDATA),
        .xillybus_S_AXI_wready(xillybus_S_AXI_WREADY),
        .xillybus_S_AXI_wstrb(xillybus_S_AXI_WSTRB),
        .xillybus_S_AXI_wvalid(xillybus_S_AXI_WVALID),
        .xillybus_bus_clk(xillybus_bus_clk),
        .xillybus_bus_rst_n(xillybus_bus_rst_n),
        .xillybus_host_interrupt(xillybus_host_interrupt), */
        
    /*    .mdio_phy_mdc(mdio_phy_mdc),
        .mdio_phy_o(mdio_phy_o),
        .mdio_phy_i(mdio_phy_i),
        .mdio_phy_t(mdio_phy_t),
        */
         .mdio_rtl_mdc(mdio_phy_mdc),
        .mdio_rtl_mdio_i(mdio_phy_i),
        .mdio_rtl_mdio_o(mdio_phy_o),
        .mdio_rtl_mdio_t(mdio_phy_t),
        .rmii2phy_txd(rmii2phy_txd),
        .rmii2phy_tx_en(rmii2phy_tx_en),
        .phy2rmii_rx_er(phy2rmii_rx_er),
        .phy2rmii_crs_dv(phy2rmii_crs_dv),
        .phy2rmii_rxd(phy2rmii_rxd),
        .ethclk50(ethclk50),
        .reset_rtl(reset_rtl)
 
        
        );
endmodule
